menosum_inst : menosum PORT MAP (
		result	 => result_sig
	);
