CONST_Value_1_inst : CONST_Value_1 PORT MAP (
		result	 => result_sig
	);
