INT31BtoFloat_inst : INT31BtoFloat PORT MAP (
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		result	 => result_sig
	);
