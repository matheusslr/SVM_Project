const_sigma_inst : const_sigma PORT MAP (
		result	 => result_sig
	);
