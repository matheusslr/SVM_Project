Convert_INT_Float_inst : Convert_INT_Float PORT MAP (
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		result	 => result_sig
	);
